module half_adder(sum,carry,a,b);
input a,b;
output sum,carry;
xor2 g1(a,b,sum);
and g2(carry,a,b);
endmodule
