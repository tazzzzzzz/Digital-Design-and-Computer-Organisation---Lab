//Module full adder.



// Module 4-bit ripple carry adder.


module fa4 (input wire [3:0] a, b, input wire cin, output wire [3:0] sum, output wire cout);

 
  // Instantiate full adder modules here.


endmodule 


    